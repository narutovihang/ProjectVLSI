*** SPICE deck for cell column4_4{lay} from library SRAM_8x8
*** Created on Sat Mar 21, 2015 16:10:37
*** Last revised on Fri Apr 03, 2015 11:32:08
*** Written on Fri Apr 03, 2015 11:32:46 by Electric VLSI Design System, 
*** version 9.05
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SRAM_8x8__NAND3 FROM CELL NAND3{lay}
.SUBCKT SRAM_8x8__NAND3 A ABC B C gnd vdd
Mncc@2 net@3 A ABC gnd NMOS L=0.6U W=3U AS=8.213P AD=2.7P PS=10.05U PD=4.8U
Mnmos@0 net@4 B net@3 gnd NMOS L=0.6U W=3U AS=2.7P AD=2.7P PS=4.8U PD=4.8U
Mnmos@2 gnd C net@4 gnd NMOS L=0.6U W=3U AS=2.7P AD=25.2P PS=4.8U PD=37.8U
Mpmos@0 ABC A vdd vdd PMOS L=0.6U W=4.5U AS=14.55P AD=8.213P PS=18.8U 
+PD=10.05U
Mpmos@1 vdd B ABC vdd PMOS L=0.6U W=4.5U AS=8.213P AD=14.55P PS=10.05U 
+PD=18.8U
Mpmos@2 ABC C vdd vdd PMOS L=0.6U W=4.5U AS=14.55P AD=8.213P PS=18.8U 
+PD=10.05U
.ENDS SRAM_8x8__NAND3

*** SUBCIRCUIT inverter1__inv FROM CELL inverter1:inv{lay}
.SUBCKT inverter1__inv gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U AS=10.35P AD=6.75P PS=18.9U PD=12.6U
Mpmos@0 out in vdd vdd PMOS L=0.6U W=6U AS=12.6P AD=6.75P PS=24.6U PD=12.6U
.ENDS inverter1__inv

*** SUBCIRCUIT SRAM_8x8__decoder_2 FROM CELL decoder_2{lay}
.SUBCKT SRAM_8x8__decoder_2 A B C Den gnd I0 I1 I2 I3 I4 I5 I6 I7 vdd
XNAND3@0 net@721 I0 net@724 net@727 gnd vdd SRAM_8x8__NAND3
XNAND3@1 net@721 I1 net@724 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@2 net@721 I2 net@5 net@727 gnd vdd SRAM_8x8__NAND3
XNAND3@3 net@721 I3 net@5 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@5 net@1 I4 net@724 net@727 gnd vdd SRAM_8x8__NAND3
XNAND3@6 net@1 I5 net@724 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@7 net@1 I6 net@5 net@727 gnd vdd SRAM_8x8__NAND3
XNAND3@8 net@1 I7 net@5 net@10 gnd vdd SRAM_8x8__NAND3
Xinv@0 gnd Den net@22 vdd inverter1__inv
Xinv@1 gnd net@1 net@721 vdd inverter1__inv
Xinv@2 gnd net@5 net@724 vdd inverter1__inv
Xinv@3 gnd net@10 net@727 vdd inverter1__inv
Mnmos@0 A Den net@1 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U PD=15.6U
Mnmos@1 B Den net@5 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U PD=15.6U
Mnmos@2 C Den net@10 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@0 A net@22 net@1 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@1 B net@22 net@5 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@2 C net@22 net@10 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
.ENDS SRAM_8x8__decoder_2

*** SUBCIRCUIT inverter1__inv_2 FROM CELL inverter1:inv_2{lay}
.SUBCKT inverter1__inv_2 gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U AS=10.35P AD=6.75P PS=18.9U PD=12.6U
Mpmos@0 out in vdd vdd PMOS L=0.6U W=6U AS=12.6P AD=6.75P PS=24.6U PD=12.6U
.ENDS inverter1__inv_2

*** TOP LEVEL CELL: column4_4{lay}
Xdecoder_@0 A B C DEN gnd net@4666 net@4673 net@4686 net@4676 net@4678 
+net@4681 net@4682 net@6205 vdd SRAM_8x8__decoder_2
Xinv_2@0 gnd net@4666 net@387 vdd inverter1__inv_2
Xinv_2@1 gnd net@4673 net@1411 vdd inverter1__inv_2
Xinv_2@2 gnd net@4686 net@1997 vdd inverter1__inv_2
Xinv_2@3 gnd net@4676 net@1803 vdd inverter1__inv_2
Xinv_2@4 gnd net@4678 net@2586 vdd inverter1__inv_2
Xinv_2@5 gnd net@4681 net@2604 vdd inverter1__inv_2
Xinv_2@6 gnd net@4682 net@3190 vdd inverter1__inv_2
Xinv_2@7 gnd net@6205 net@2996 vdd inverter1__inv_2
Mnmos@18 gnd net@339 net@329 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@19 gnd net@329 net@339 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@20 net@480 net@387 net@329 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@21 net@481 net@387 net@339 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@22 gnd net@586 net@584 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@23 gnd net@584 net@586 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@24 net@613 net@387 net@584 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@25 net@614 net@387 net@586 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=73.064P 
+PS=16.05U PD=57.436U
Mnmos@26 gnd net@634 net@632 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@27 gnd net@632 net@634 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@28 net@661 net@387 net@632 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@29 net@662 net@387 net@634 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@30 gnd net@683 net@681 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@31 gnd net@681 net@683 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@32 net@710 net@387 net@681 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@33 net@711 net@387 net@683 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@34 gnd net@727 net@725 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@35 gnd net@725 net@727 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@36 net@754 net@387 net@725 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@37 net@755 net@387 net@727 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@38 gnd net@771 net@769 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@39 gnd net@769 net@771 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@40 net@798 net@387 net@769 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@41 net@799 net@387 net@771 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@50 gnd net@924 net@922 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@51 gnd net@922 net@924 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@52 net@951 net@387 net@922 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@53 net@952 net@387 net@924 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@54 gnd net@971 net@969 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@55 gnd net@969 net@971 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@56 net@998 net@387 net@969 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@57 net@999 net@387 net@971 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@90 gnd net@1415 net@1413 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@91 gnd net@1413 net@1415 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@92 net@480 net@1411 net@1413 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@93 net@481 net@1411 net@1415 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@94 gnd net@1458 net@1456 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@95 gnd net@1456 net@1458 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@96 net@613 net@1411 net@1456 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@97 net@614 net@1411 net@1458 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=73.064P PS=16.05U PD=57.436U
Mnmos@98 gnd net@1504 net@1502 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@99 gnd net@1502 net@1504 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@100 net@661 net@1411 net@1502 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@101 net@662 net@1411 net@1504 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@102 gnd net@1549 net@1547 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@103 gnd net@1547 net@1549 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@104 net@710 net@1411 net@1547 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@105 net@711 net@1411 net@1549 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@106 gnd net@1593 net@1591 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@107 gnd net@1591 net@1593 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@108 net@754 net@1411 net@1591 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@109 net@755 net@1411 net@1593 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@110 gnd net@1637 net@1635 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@111 gnd net@1635 net@1637 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@112 net@798 net@1411 net@1635 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@113 net@799 net@1411 net@1637 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@114 gnd net@1693 net@1691 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@115 gnd net@1691 net@1693 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@116 net@951 net@1411 net@1691 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@117 net@952 net@1411 net@1693 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@118 gnd net@1400 net@1403 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@119 gnd net@1403 net@1400 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@120 net@998 net@1411 net@1403 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@121 net@999 net@1411 net@1400 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@122 gnd net@1987 net@1985 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@123 gnd net@1985 net@1987 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@124 net@480 net@1997 net@1985 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@125 net@481 net@1997 net@1987 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@126 gnd net@2030 net@2028 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@127 gnd net@2028 net@2030 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@128 net@613 net@1997 net@2028 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@129 net@614 net@1997 net@2030 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=73.064P PS=16.05U PD=57.436U
Mnmos@130 gnd net@2076 net@2074 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@131 gnd net@2074 net@2076 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@132 net@661 net@1997 net@2074 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@133 net@662 net@1997 net@2076 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@134 gnd net@2121 net@2119 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@135 gnd net@2119 net@2121 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@136 net@710 net@1997 net@2119 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@137 net@711 net@1997 net@2121 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@138 gnd net@2165 net@2163 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@139 gnd net@2163 net@2165 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@140 net@754 net@1997 net@2163 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@141 net@755 net@1997 net@2165 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@142 gnd net@2209 net@2207 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@143 gnd net@2207 net@2209 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@144 net@798 net@1997 net@2207 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@145 net@799 net@1997 net@2209 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@146 gnd net@2265 net@2263 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@147 gnd net@2263 net@2265 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@148 net@951 net@1997 net@2263 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@149 net@952 net@1997 net@2265 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@150 gnd net@2312 net@2310 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@151 gnd net@2310 net@2312 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@152 net@998 net@1997 net@2310 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@153 net@999 net@1997 net@2312 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@154 gnd net@2379 net@2377 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@155 gnd net@2377 net@2379 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@156 net@480 net@1803 net@2377 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@157 net@481 net@1803 net@2379 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@158 gnd net@2422 net@2420 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@159 gnd net@2420 net@2422 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@160 net@613 net@1803 net@2420 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@161 net@614 net@1803 net@2422 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=73.064P PS=16.05U PD=57.436U
Mnmos@162 gnd net@2468 net@2466 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@163 gnd net@2466 net@2468 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@164 net@661 net@1803 net@2466 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@165 net@662 net@1803 net@2468 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@166 gnd net@1785 net@1786 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@167 gnd net@1786 net@1785 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@168 net@710 net@1803 net@1786 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@169 net@711 net@1803 net@1785 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@170 gnd net@1793 net@1791 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@171 gnd net@1791 net@1793 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@172 net@754 net@1803 net@1791 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@173 net@755 net@1803 net@1793 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@174 gnd net@1837 net@1835 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@175 gnd net@1835 net@1837 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@176 net@798 net@1803 net@1835 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@177 net@799 net@1803 net@1837 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@178 gnd net@1893 net@1891 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@179 gnd net@1891 net@1893 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@180 net@951 net@1803 net@1891 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@181 net@952 net@1803 net@1893 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@182 gnd net@1940 net@1938 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@183 gnd net@1938 net@1940 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@184 net@998 net@1803 net@1938 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@185 net@999 net@1803 net@1940 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@186 gnd p47 o47 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@187 gnd o47 p47 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@188 net@480 net@2586 o47 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@189 net@481 net@2586 p47 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@190 gnd p46 net@3802 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@191 gnd net@3802 p46 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@192 net@613 net@2586 net@3802 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@193 net@614 net@2586 p46 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=73.064P 
+PS=16.05U PD=57.436U
Mnmos@194 gnd p45 net@3848 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@195 gnd net@3848 p45 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@196 net@661 net@2586 net@3848 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@197 net@662 net@2586 p45 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@198 gnd p44 net@3893 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@199 gnd net@3893 p44 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@200 net@710 net@2586 net@3893 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@201 net@711 net@2586 p44 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@202 gnd p43 net@3937 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@203 gnd net@3937 p43 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@204 net@754 net@2586 net@3937 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@205 net@755 net@2586 p43 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@206 gnd p42 net@3981 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@207 gnd net@3981 p42 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@208 net@798 net@2586 net@3981 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@209 net@799 net@2586 p42 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@210 gnd p41 net@4037 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@211 gnd net@4037 p41 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@212 net@951 net@2586 net@4037 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@213 net@952 net@2586 p41 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@214 gnd p40 o40 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@215 gnd o40 p40 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@216 net@998 net@2586 o40 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@217 net@999 net@2586 p40 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@218 gnd p57 o57 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@219 gnd o57 p57 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@220 net@480 net@2604 o57 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@221 net@481 net@2604 p57 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@222 gnd p56 net@2649 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@223 gnd net@2649 p56 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@224 net@613 net@2604 net@2649 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@225 net@614 net@2604 p56 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=73.064P 
+PS=16.05U PD=57.436U
Mnmos@226 gnd p55 net@2695 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@227 gnd net@2695 p55 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@228 net@661 net@2604 net@2695 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@229 net@662 net@2604 p55 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@230 gnd p54 net@2740 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@231 gnd net@2740 p54 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@232 net@710 net@2604 net@2740 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@233 net@711 net@2604 p54 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@234 gnd p53 net@2784 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@235 gnd net@2784 p53 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@236 net@754 net@2604 net@2784 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@237 net@755 net@2604 p53 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@238 gnd p52 net@2828 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@239 gnd net@2828 p52 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@240 net@798 net@2604 net@2828 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@241 net@799 net@2604 p52 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@242 gnd p51 net@2884 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@243 gnd net@2884 p51 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@244 net@951 net@2604 net@2884 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@245 net@952 net@2604 p51 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@246 gnd p50 o50 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@247 gnd o50 p50 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@248 net@998 net@2604 o50 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@249 net@999 net@2604 p50 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@250 gnd net@3180 net@3178 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@251 gnd net@3178 net@3180 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@252 net@480 net@3190 net@3178 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@253 net@481 net@3190 net@3180 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@254 gnd net@3223 net@3221 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@255 gnd net@3221 net@3223 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@256 net@613 net@3190 net@3221 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@257 net@614 net@3190 net@3223 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=73.064P PS=16.05U PD=57.436U
Mnmos@258 gnd net@3269 net@3267 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@259 gnd net@3267 net@3269 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@260 net@661 net@3190 net@3267 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@261 net@662 net@3190 net@3269 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@262 gnd net@3314 net@3312 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@263 gnd net@3312 net@3314 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@264 net@710 net@3190 net@3312 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@265 net@711 net@3190 net@3314 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@266 gnd net@3358 net@3356 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@267 gnd net@3356 net@3358 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@268 net@754 net@3190 net@3356 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@269 net@755 net@3190 net@3358 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@270 gnd net@3402 net@3400 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@271 gnd net@3400 net@3402 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@272 net@798 net@3190 net@3400 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@273 net@799 net@3190 net@3402 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@274 gnd net@3458 net@3456 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@275 gnd net@3456 net@3458 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@276 net@951 net@3190 net@3456 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@277 net@952 net@3190 net@3458 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@278 gnd net@3505 net@3503 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@279 gnd net@3503 net@3505 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@280 net@998 net@3190 net@3503 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@281 net@999 net@3190 net@3505 gnd NMOS L=0.6U W=4.5U AS=8.287P 
+AD=32.973P PS=16.05U PD=30.164U
Mnmos@282 gnd p77 o77 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@283 gnd o77 p77 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@284 net@480 net@2996 o77 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@285 net@481 net@2996 p77 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@286 gnd p76 net@3613 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@287 gnd net@3613 p76 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@288 net@613 net@2996 net@3613 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@289 net@614 net@2996 p76 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=73.064P 
+PS=16.05U PD=57.436U
Mnmos@290 gnd p75 net@3659 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@291 gnd net@3659 p75 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@292 net@661 net@2996 net@3659 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@293 net@662 net@2996 p75 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@294 gnd p74 net@2979 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@295 gnd net@2979 p74 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@296 net@710 net@2996 net@2979 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@297 net@711 net@2996 p74 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@298 gnd p73 net@2984 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@299 gnd net@2984 p73 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@300 net@754 net@2996 net@2984 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@301 net@755 net@2996 p73 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@302 gnd p72 net@3028 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@303 gnd net@3028 p72 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@304 net@798 net@2996 net@3028 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@305 net@799 net@2996 p72 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@306 gnd p71 net@3084 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P 
+PS=16.45U PD=42.077U
Mnmos@307 gnd net@3084 p71 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P 
+PS=16.05U PD=42.077U
Mnmos@308 net@951 net@2996 net@3084 gnd NMOS L=0.6U W=4.5U AS=9.037P 
+AD=32.973P PS=16.45U PD=30.164U
Mnmos@309 net@952 net@2996 p71 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@310 gnd p70 o70 gnd NMOS L=0.6U W=11.25U AS=9.037P AD=28.36P PS=16.45U 
+PD=42.077U
Mnmos@311 gnd o70 p70 gnd NMOS L=0.6U W=11.25U AS=8.287P AD=28.36P PS=16.05U 
+PD=42.077U
Mnmos@312 net@998 net@2996 o70 gnd NMOS L=0.6U W=4.5U AS=9.037P AD=32.973P 
+PS=16.45U PD=30.164U
Mnmos@313 net@999 net@2996 p70 gnd NMOS L=0.6U W=4.5U AS=8.287P AD=32.973P 
+PS=16.05U PD=30.164U
Mnmos@314 net@6542 qo net@7169 gnd NMOS L=0.6U W=3U AS=5.362P AD=64.575P 
+PS=11.35U PD=75.45U
Mnmos@315 qo net@6542 net@7169 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.787P 
+PS=11.35U PD=74.55U
Mnmos@316 gnd SAE net@7169 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@317 net@7127 WE net@6542 gnd NMOS L=0.6U W=67.5U AS=64.575P AD=61.155P 
+PS=75.45U PD=136.8U
Mnmos@318 gnd d0 net@7127 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@319 net@7132 WE qo gnd NMOS L=0.6U W=67.5U AS=63.787P AD=61.222P 
+PS=74.55U PD=136.95U
Mnmos@320 gnd net@7143 net@7132 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@321 gnd d0 net@7143 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@322 net@7227 q1 net@7279 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.675P 
+PS=11.35U PD=74.25U
Mnmos@323 q1 net@7227 net@7279 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.45P 
+PS=11.35U PD=74.1U
Mnmos@324 gnd SAE net@7279 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@325 net@7234 WE net@7227 gnd NMOS L=0.6U W=67.5U AS=63.675P AD=61.155P 
+PS=74.25U PD=136.8U
Mnmos@326 gnd d1 net@7234 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@327 net@7240 WE q1 gnd NMOS L=0.6U W=67.5U AS=63.45P AD=61.222P 
+PS=74.1U PD=136.95U
Mnmos@328 gnd net@7251 net@7240 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@329 gnd d1 net@7251 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@330 net@6414 q2 net@6837 gnd NMOS L=0.6U W=3U AS=5.362P AD=64.575P 
+PS=11.35U PD=75.45U
Mnmos@331 q2 net@6414 net@6837 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.787P 
+PS=11.35U PD=74.55U
Mnmos@332 gnd SAE net@6837 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@333 net@7081 WE net@6414 gnd NMOS L=0.6U W=67.5U AS=64.575P AD=61.155P 
+PS=75.45U PD=136.8U
Mnmos@334 gnd d2 net@7081 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@335 net@6438 WE q2 gnd NMOS L=0.6U W=67.5U AS=63.787P AD=61.222P 
+PS=74.55U PD=136.95U
Mnmos@336 gnd net@6549 net@6438 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@337 gnd d2 net@6549 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@338 net@6419 q3 net@6468 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.675P 
+PS=11.35U PD=74.25U
Mnmos@339 q3 net@6419 net@6468 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.45P 
+PS=11.35U PD=74.1U
Mnmos@340 gnd SAE net@6468 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@341 net@6423 WE net@6419 gnd NMOS L=0.6U W=67.5U AS=63.675P AD=61.155P 
+PS=74.25U PD=136.8U
Mnmos@342 gnd d3 net@6423 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@343 net@6429 WE q3 gnd NMOS L=0.6U W=67.5U AS=63.45P AD=61.222P 
+PS=74.1U PD=136.95U
Mnmos@344 gnd net@6440 net@6429 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@345 gnd d3 net@6440 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@346 net@6769 q4 net@6822 gnd NMOS L=0.6U W=3U AS=5.362P AD=64.575P 
+PS=11.35U PD=75.45U
Mnmos@347 q4 net@6769 net@6822 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.787P 
+PS=11.35U PD=74.55U
Mnmos@348 gnd SAE net@6822 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@349 net@6777 WE net@6769 gnd NMOS L=0.6U W=67.5U AS=64.575P AD=61.155P 
+PS=75.45U PD=136.8U
Mnmos@350 gnd d4 net@6777 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@351 net@6783 WE q4 gnd NMOS L=0.6U W=67.5U AS=63.787P AD=61.222P 
+PS=74.55U PD=136.95U
Mnmos@352 gnd net@6794 net@6783 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@353 gnd d4 net@6794 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@354 net@6879 q5 net@6932 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.675P 
+PS=11.35U PD=74.25U
Mnmos@355 q5 net@6879 net@6932 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.45P 
+PS=11.35U PD=74.1U
Mnmos@356 gnd SAE net@6932 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@357 net@6887 WE net@6879 gnd NMOS L=0.6U W=67.5U AS=63.675P AD=61.155P 
+PS=74.25U PD=136.8U
Mnmos@358 gnd d5 net@6887 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@359 net@6892 WE q5 gnd NMOS L=0.6U W=67.5U AS=63.45P AD=61.222P 
+PS=74.1U PD=136.95U
Mnmos@360 gnd net@6903 net@6892 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@361 gnd d5 net@6903 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@362 net@6536 q6 net@6590 gnd NMOS L=0.6U W=3U AS=5.362P AD=64.575P 
+PS=11.35U PD=75.45U
Mnmos@363 q6 net@6536 net@6590 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.81P 
+PS=11.35U PD=74.625U
Mnmos@364 gnd SAE net@6590 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@365 net@6545 WE net@6536 gnd NMOS L=0.6U W=67.5U AS=64.575P AD=61.155P 
+PS=75.45U PD=136.8U
Mnmos@366 gnd d6 net@6545 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@367 net@6551 WE q6 gnd NMOS L=0.6U W=67.5U AS=63.81P AD=61.222P 
+PS=74.625U PD=136.95U
Mnmos@368 gnd net@6562 net@6551 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@369 gnd d6 net@6562 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mnmos@370 net@6648 q7 net@6702 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.675P 
+PS=11.35U PD=74.25U
Mnmos@371 q7 net@6648 net@6702 gnd NMOS L=0.6U W=3U AS=5.362P AD=63.45P 
+PS=11.35U PD=74.1U
Mnmos@372 gnd SAE net@6702 gnd NMOS L=0.6U W=3U AS=5.362P AD=28.36P PS=11.35U 
+PD=42.077U
Mnmos@373 net@6656 WE net@6648 gnd NMOS L=0.6U W=67.5U AS=63.675P AD=61.155P 
+PS=74.25U PD=136.8U
Mnmos@374 gnd d7 net@6656 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=28.36P 
+PS=136.8U PD=42.077U
Mnmos@375 net@6663 WE q7 gnd NMOS L=0.6U W=67.5U AS=63.45P AD=61.222P 
+PS=74.1U PD=136.95U
Mnmos@376 gnd net@6674 net@6663 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=28.36P 
+PS=136.95U PD=42.077U
Mnmos@377 gnd d7 net@6674 gnd NMOS L=0.6U W=3U AS=10.125P AD=28.36P PS=14.1U 
+PD=42.077U
Mpmos@10 net@329 net@339 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@11 vdd net@329 net@339 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@12 net@584 net@586 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@13 vdd net@584 net@586 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@14 net@632 net@634 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@15 vdd net@632 net@634 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@16 net@681 net@683 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@17 vdd net@681 net@683 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@18 net@725 net@727 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@19 vdd net@725 net@727 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@20 net@769 net@771 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@21 vdd net@769 net@771 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@26 net@922 net@924 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@27 vdd net@922 net@924 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@28 net@969 net@971 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@29 vdd net@969 net@971 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@46 net@1413 net@1415 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@47 vdd net@1413 net@1415 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@48 net@1456 net@1458 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@49 vdd net@1456 net@1458 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@50 net@1502 net@1504 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@51 vdd net@1502 net@1504 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@52 net@1547 net@1549 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@53 vdd net@1547 net@1549 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@54 net@1591 net@1593 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@55 vdd net@1591 net@1593 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@56 net@1635 net@1637 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@57 vdd net@1635 net@1637 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@58 net@1691 net@1693 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@59 vdd net@1691 net@1693 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@60 net@1403 net@1400 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@61 vdd net@1403 net@1400 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@62 net@1985 net@1987 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@63 vdd net@1985 net@1987 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@64 net@2028 net@2030 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@65 vdd net@2028 net@2030 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@66 net@2074 net@2076 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@67 vdd net@2074 net@2076 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@68 net@2119 net@2121 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@69 vdd net@2119 net@2121 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@70 net@2163 net@2165 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@71 vdd net@2163 net@2165 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@72 net@2207 net@2209 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@73 vdd net@2207 net@2209 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@74 net@2263 net@2265 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@75 vdd net@2263 net@2265 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@76 net@2310 net@2312 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@77 vdd net@2310 net@2312 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@78 net@2377 net@2379 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@79 vdd net@2377 net@2379 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@80 net@2420 net@2422 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@81 vdd net@2420 net@2422 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@82 net@2466 net@2468 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@83 vdd net@2466 net@2468 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@84 net@1786 net@1785 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@85 vdd net@1786 net@1785 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@86 net@1791 net@1793 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@87 vdd net@1791 net@1793 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@88 net@1835 net@1837 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@89 vdd net@1835 net@1837 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@90 net@1891 net@1893 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@91 vdd net@1891 net@1893 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@92 net@1938 net@1940 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@93 vdd net@1938 net@1940 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@94 o47 p47 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@95 vdd o47 p47 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@96 net@3802 p46 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@97 vdd net@3802 p46 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@98 net@3848 p45 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@99 vdd net@3848 p45 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@100 net@3893 p44 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@101 vdd net@3893 p44 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@102 net@3937 p43 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@103 vdd net@3937 p43 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@104 net@3981 p42 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@105 vdd net@3981 p42 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@106 net@4037 p41 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@107 vdd net@4037 p41 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@108 o40 p40 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@109 vdd o40 p40 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@110 o57 p57 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@111 vdd o57 p57 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@112 net@2649 p56 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@113 vdd net@2649 p56 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@114 net@2695 p55 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@115 vdd net@2695 p55 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@116 net@2740 p54 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@117 vdd net@2740 p54 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@118 net@2784 p53 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@119 vdd net@2784 p53 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@120 net@2828 p52 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@121 vdd net@2828 p52 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@122 net@2884 p51 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@123 vdd net@2884 p51 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@124 o50 p50 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@125 vdd o50 p50 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@126 net@3178 net@3180 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@127 vdd net@3178 net@3180 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@128 net@3221 net@3223 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@129 vdd net@3221 net@3223 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@130 net@3267 net@3269 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@131 vdd net@3267 net@3269 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@132 net@3312 net@3314 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@133 vdd net@3312 net@3314 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@134 net@3356 net@3358 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@135 vdd net@3356 net@3358 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@136 net@3400 net@3402 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@137 vdd net@3400 net@3402 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@138 net@3456 net@3458 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@139 vdd net@3456 net@3458 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@140 net@3503 net@3505 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@141 vdd net@3503 net@3505 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@142 o77 p77 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@143 vdd o77 p77 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@144 net@3613 p76 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@145 vdd net@3613 p76 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@146 net@3659 p75 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@147 vdd net@3659 p75 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@148 net@2979 p74 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@149 vdd net@2979 p74 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@150 net@2984 p73 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@151 vdd net@2984 p73 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@152 net@3028 p72 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@153 vdd net@3028 p72 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@154 net@3084 p71 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P 
+PS=31.257U PD=16.45U
Mpmos@155 vdd net@3084 p71 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P 
+PS=16.05U PD=31.257U
Mpmos@156 o70 p70 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=9.037P PS=31.257U 
+PD=16.45U
Mpmos@157 vdd o70 p70 vdd PMOS L=0.6U W=3U AS=8.287P AD=24.117P PS=16.05U 
+PD=31.257U
Mpmos@198 vdd P net@999 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@199 net@998 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@200 net@999 P net@998 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@201 vdd P net@952 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@202 net@951 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@203 net@952 P net@951 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@207 vdd P net@755 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@208 net@754 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@209 net@755 P net@754 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@210 vdd P net@711 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@211 net@710 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@212 net@711 P net@710 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@213 vdd P net@662 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@214 net@661 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@215 net@662 P net@661 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@216 vdd P net@481 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@217 net@480 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@218 net@481 P net@480 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U
Mpmos@219 vdd P net@614 vdd PMOS L=0.6U W=42U AS=73.064P AD=24.117P 
+PS=57.436U PD=31.257U
Mpmos@220 net@613 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@221 net@614 P net@613 vdd PMOS L=0.6U W=42U AS=32.973P AD=73.064P 
+PS=30.164U PD=57.436U
Mpmos@222 net@6542 qo vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=64.575P 
+PS=31.257U PD=75.45U
Mpmos@223 qo net@6542 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.787P 
+PS=31.257U PD=74.55U
Mpmos@224 net@6542 SAE net@999 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=64.575P 
+PS=30.164U PD=75.45U
Mpmos@225 qo SAE net@998 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.787P 
+PS=30.164U PD=74.55U
Mpmos@226 vdd d0 net@7143 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@227 net@7227 q1 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.675P 
+PS=31.257U PD=74.25U
Mpmos@228 q1 net@7227 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.45P 
+PS=31.257U PD=74.1U
Mpmos@229 net@7227 SAE net@952 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.675P 
+PS=30.164U PD=74.25U
Mpmos@230 q1 SAE net@951 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.45P 
+PS=30.164U PD=74.1U
Mpmos@231 vdd d1 net@7251 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@232 net@6414 q2 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=64.575P 
+PS=31.257U PD=75.45U
Mpmos@233 q2 net@6414 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.787P 
+PS=31.257U PD=74.55U
Mpmos@234 net@6414 SAE net@799 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=64.575P 
+PS=30.164U PD=75.45U
Mpmos@235 q2 SAE net@798 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.787P 
+PS=30.164U PD=74.55U
Mpmos@236 vdd d2 net@6549 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@237 net@6419 q3 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.675P 
+PS=31.257U PD=74.25U
Mpmos@238 q3 net@6419 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.45P 
+PS=31.257U PD=74.1U
Mpmos@239 net@6419 SAE net@755 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.675P 
+PS=30.164U PD=74.25U
Mpmos@240 q3 SAE net@754 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.45P 
+PS=30.164U PD=74.1U
Mpmos@241 vdd d3 net@6440 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@242 net@6769 q4 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=64.575P 
+PS=31.257U PD=75.45U
Mpmos@243 q4 net@6769 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.787P 
+PS=31.257U PD=74.55U
Mpmos@244 net@6769 SAE net@711 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=64.575P 
+PS=30.164U PD=75.45U
Mpmos@245 q4 SAE net@710 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.787P 
+PS=30.164U PD=74.55U
Mpmos@246 vdd d4 net@6794 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@247 net@6879 q5 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.675P 
+PS=31.257U PD=74.25U
Mpmos@248 q5 net@6879 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.45P 
+PS=31.257U PD=74.1U
Mpmos@249 net@6879 SAE net@662 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.675P 
+PS=30.164U PD=74.25U
Mpmos@250 q5 SAE net@661 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.45P 
+PS=30.164U PD=74.1U
Mpmos@251 vdd d5 net@6903 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@252 net@6536 q6 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=64.575P 
+PS=31.257U PD=75.45U
Mpmos@253 q6 net@6536 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.81P 
+PS=31.257U PD=74.625U
Mpmos@254 net@6536 SAE net@614 vdd PMOS L=0.6U W=67.5U AS=73.064P AD=64.575P 
+PS=57.436U PD=75.45U
Mpmos@255 q6 SAE net@613 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.81P 
+PS=30.164U PD=74.625U
Mpmos@256 vdd d6 net@6562 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@257 net@6648 q7 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.675P 
+PS=31.257U PD=74.25U
Mpmos@258 q7 net@6648 vdd vdd PMOS L=0.6U W=3U AS=24.117P AD=63.45P 
+PS=31.257U PD=74.1U
Mpmos@259 net@6648 SAE net@481 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.675P 
+PS=30.164U PD=74.25U
Mpmos@260 q7 SAE net@480 vdd PMOS L=0.6U W=67.5U AS=32.973P AD=63.45P 
+PS=30.164U PD=74.1U
Mpmos@261 vdd d7 net@6674 vdd PMOS L=0.6U W=6U AS=10.125P AD=24.117P PS=14.1U 
+PD=31.257U
Mpmos@262 vdd P net@799 vdd PMOS L=0.6U W=42U AS=32.973P AD=24.117P 
+PS=30.164U PD=31.257U
Mpmos@263 net@798 P vdd vdd PMOS L=0.6U W=42U AS=24.117P AD=32.973P 
+PS=31.257U PD=30.164U
Mpmos@264 net@799 P net@798 vdd PMOS L=0.6U W=42U AS=32.973P AD=32.973P 
+PS=30.164U PD=30.164U

* Spice Code nodes in cell cell 'column4_4{lay}'
vdd vdd 0 dc 5
va A 0 DC 0 pwl 100n 0 110n 5 150n 5 160n 0 200n 0 210n 5
vb B 0 DC 0 pwl 100n 5 110n 0 200n 0 210n 5 350n 5 360n 0 500n 0 510n 5
vc C 0 DC 0 pwl 100n 0 110n 5 350n 5 360n 0 500n 0 510n 5
vp P 0 DC 0 pwl 50n 5 60n 0 100n 0 110n 5 200n 5 210n 0 250n 0 260n 5 350n 5 
+360n 0 400n 0 410n 5 500n 5 510n 0 550n 0 560n 5
vwe WE 0 DC 0 pwl 100n 5 110n 0 250n 0 260n 5 300n 5 310n 0
vsae SAE 0 DC 0 pwl 100n 5 110n 0 150n 0 160n 5 250n 5 260n 0 300n 0 310n 5 
+400n 5 410n 0 450n 0 460n 5 550n 5 560n 0 600n 0 610n 5
vden DEN 0 dc 0 pwl 100n 0 110n 5 150n 5 160n 0 250n 0 260n 5 300n 5 310n 0 
+400n 0 410n 5 450n 5 460n 0 550n 0 560n 5 600n 5 610n 0
vd0 d0 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd1 d1 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd2 d2 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd3 d3 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd4 d4 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd5 d5 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd6 d6 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd7 d7 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
.IC V(p50)=0 V(p51)=0 V(p52)=0 V(p53)=0 V(p54)=0 V(p55)=0 V(p56)=0 V(p57)=0 
+V(p40)=0 V(p41)=0 V(p42)=0 V(p43)=0 V(p44)=0 V(p45)=0 V(p46)=0 V(p47)=0 
+V(p70)=0 V(p71)=0 V(p72)=0 V(p73)=0 V(p74)=0 V(p75)=0 V(p76)=0 V(p77)=0
.tran 0 800ns
.include C5_models.txt
.END
