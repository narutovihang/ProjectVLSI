*** SPICE deck for cell decoder{sch} from library SRAM_8x8
*** Created on Tue Dec 30, 2014 13:22:16
*** Last revised on Wed Mar 25, 2015 15:26:48
*** Written on Wed Mar 25, 2015 15:26:51 by Electric VLSI Design System, 
*** version 9.05
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SRAM_8x8__NAND3 FROM CELL NAND3{sch}
.SUBCKT SRAM_8x8__NAND3 A ABC B C
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 ABC A net@40 gnd NMOS L=0.4U W=2U
Mnmos@1 net@40 B net@43 gnd NMOS L=0.4U W=2U
Mnmos@2 net@43 C gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd A ABC vdd PMOS L=0.4U W=3U
Mpmos@1 vdd B ABC vdd PMOS L=0.4U W=3U
Mpmos@2 vdd C ABC vdd PMOS L=0.4U W=3U
.ENDS SRAM_8x8__NAND3

*** SUBCIRCUIT SRAM_8x8__inv FROM CELL inv{sch}
.SUBCKT SRAM_8x8__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=4U
.ENDS SRAM_8x8__inv

.global gnd vdd

*** TOP LEVEL CELL: decoder{sch}
Mnmos@0 net@40 Den A gnd NMOS L=0.4U W=0.4U
Mnmos@1 net@38 Den B gnd NMOS L=0.4U W=0.4U
Mnmos@2 net@36 Den C gnd NMOS L=0.4U W=0.4U
Mpmos@0 A net@166 net@40 vdd PMOS L=0.4U W=0.4U
Mpmos@1 B net@166 net@38 vdd PMOS L=0.4U W=0.4U
Mpmos@2 C net@166 net@36 vdd PMOS L=0.4U W=0.4U
XNAND3@0 net@40 I7 net@38 net@36 SRAM_8x8__NAND3
XNAND3@1 net@40 I6 net@38 net@94 SRAM_8x8__NAND3
XNAND3@2 net@40 I5 net@53 net@36 SRAM_8x8__NAND3
XNAND3@3 net@40 I4 net@53 net@94 SRAM_8x8__NAND3
XNAND3@4 net@184 I3 net@38 net@36 SRAM_8x8__NAND3
XNAND3@5 net@184 I2 net@38 net@94 SRAM_8x8__NAND3
XNAND3@6 net@184 I1 net@53 net@36 SRAM_8x8__NAND3
XNAND3@7 net@184 I0 net@53 net@94 SRAM_8x8__NAND3
Xinv@5 net@40 net@184 SRAM_8x8__inv
Xinv@6 net@38 net@53 SRAM_8x8__inv
Xinv@7 net@36 net@94 SRAM_8x8__inv
Xinv@8 Den net@166 SRAM_8x8__inv

* Spice Code nodes in cell cell 'decoder{sch}'
vdd vdd 0 dc 5
v1 A 0 dc 0
v2 B 0 dc 0
v3 C 0 dc 5
.tran 800ns
.include C5_models.txt
.END
