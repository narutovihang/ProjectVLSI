*** SPICE deck for cell column4{lay} from library SRAM_8x8
*** Created on Tue Mar 24, 2015 17:42:07
*** Last revised on Wed Apr 01, 2015 19:53:26
*** Written on Wed Apr 01, 2015 19:55:44 by Electric VLSI Design System, 
*** version 9.05
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Cell_Copy__cell2 FROM CELL Cell_Copy:cell2{lay}
.SUBCKT Cell_Copy__cell2 B Bb gnd n q vdd W
Mnmos@0 q n gnd gnd NMOS L=0.6U W=11.25U AS=19.125P AD=10.783P PS=37.8U 
+PD=19.85U
Mnmos@1 gnd q n gnd NMOS L=0.6U W=11.25U AS=9.617P AD=19.125P PS=18.55U 
+PD=37.8U
Mnmos@4 Bb W q gnd NMOS L=0.6U W=4.5U AS=10.783P AD=8.055P PS=19.85U PD=18.9U
Mnmos@5 B W n gnd NMOS L=0.6U W=4.5U AS=9.617P AD=6.3P PS=18.55U PD=13.8U
Mpmos@0 q n vdd vdd PMOS L=0.6U W=3U AS=11.7P AD=10.783P PS=21.3U PD=19.85U
Mpmos@1 vdd q n vdd PMOS L=0.6U W=3U AS=9.617P AD=11.7P PS=18.55U PD=21.3U
.ENDS Cell_Copy__cell2

*** SUBCIRCUIT SRAM_8x8__NAND3 FROM CELL NAND3{lay}
.SUBCKT SRAM_8x8__NAND3 A ABC B C gnd vdd
Mncc@2 net@3 A ABC gnd NMOS L=0.6U W=3U AS=8.213P AD=2.7P PS=10.05U PD=4.8U
Mnmos@0 net@4 B net@3 gnd NMOS L=0.6U W=3U AS=2.7P AD=2.7P PS=4.8U PD=4.8U
Mnmos@2 gnd C net@4 gnd NMOS L=0.6U W=3U AS=2.7P AD=25.2P PS=4.8U PD=37.8U
Mpmos@0 ABC A vdd vdd PMOS L=0.6U W=4.5U AS=14.55P AD=8.213P PS=18.8U 
+PD=10.05U
Mpmos@1 vdd B ABC vdd PMOS L=0.6U W=4.5U AS=8.213P AD=14.55P PS=10.05U 
+PD=18.8U
Mpmos@2 ABC C vdd vdd PMOS L=0.6U W=4.5U AS=14.55P AD=8.213P PS=18.8U 
+PD=10.05U
.ENDS SRAM_8x8__NAND3

*** SUBCIRCUIT inverter1__inv FROM CELL inverter1:inv{lay}
.SUBCKT inverter1__inv gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U AS=10.35P AD=6.75P PS=18.9U PD=12.6U
Mpmos@0 out in vdd vdd PMOS L=0.6U W=6U AS=12.6P AD=6.75P PS=24.6U PD=12.6U
.ENDS inverter1__inv

*** SUBCIRCUIT SRAM_8x8__decoder FROM CELL decoder{lay}
.SUBCKT SRAM_8x8__decoder A B C Den gnd I0 I1 I2 I3 I4 I5 I6 I7 vdd
XNAND3@0 net@71 I0 net@88 net@99 gnd vdd SRAM_8x8__NAND3
XNAND3@1 net@71 I1 net@88 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@2 net@71 I2 net@5 net@99 gnd vdd SRAM_8x8__NAND3
XNAND3@3 net@71 I3 net@5 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@5 net@1 I4 net@88 net@99 gnd vdd SRAM_8x8__NAND3
XNAND3@6 net@1 I5 net@88 net@10 gnd vdd SRAM_8x8__NAND3
XNAND3@7 net@1 I6 net@5 net@99 gnd vdd SRAM_8x8__NAND3
XNAND3@8 net@1 I7 net@5 net@10 gnd vdd SRAM_8x8__NAND3
Xinv@0 gnd Den net@22 vdd inverter1__inv
Xinv@1 gnd net@1 net@71 vdd inverter1__inv
Xinv@2 gnd net@5 net@88 vdd inverter1__inv
Xinv@3 gnd net@10 net@99 vdd inverter1__inv
Mnmos@0 A Den net@1 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U PD=15.6U
Mnmos@1 B Den net@5 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U PD=15.6U
Mnmos@2 C Den net@10 gnd NMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@0 A net@22 net@1 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@1 B net@22 net@5 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
Mpmos@2 C net@22 net@10 vdd PMOS L=0.6U W=0.9U AS=2.52P AD=7.02P PS=6.6U 
+PD=15.6U
.ENDS SRAM_8x8__decoder

*** SUBCIRCUIT SRAM_8x8__sense_amp FROM CELL sense_amp{lay}
.SUBCKT SRAM_8x8__sense_amp B Bb D gnd Q SAE vdd WE
Mnmos@6 net@212 Q net@136 gnd NMOS L=0.6U W=3U AS=63.225P AD=7.545P PS=73.95U 
+PD=16.2U
Mnmos@7 net@212 net@136 Q gnd NMOS L=0.6U W=3U AS=63.225P AD=7.545P PS=73.95U 
+PD=16.2U
Mnmos@8 gnd SAE net@212 gnd NMOS L=0.6U W=3U AS=7.545P AD=76.388P PS=16.2U 
+PD=94.65U
Mnmos@9 gnd D net@221 gnd NMOS L=0.6U W=3U AS=7.425P AD=76.388P PS=12.3U 
+PD=94.65U
Mnmos@12 net@275 WE net@136 gnd NMOS L=0.6U W=67.5U AS=63.225P AD=61.155P 
+PS=73.95U PD=136.8U
Mnmos@13 gnd D net@275 gnd NMOS L=0.6U W=67.5U AS=61.155P AD=76.388P 
+PS=136.8U PD=94.65U
Mnmos@14 net@281 WE Q gnd NMOS L=0.6U W=67.5U AS=63.225P AD=61.222P PS=73.95U 
+PD=136.95U
Mnmos@15 gnd net@221 net@281 gnd NMOS L=0.6U W=67.5U AS=61.222P AD=76.388P 
+PS=136.95U PD=94.65U
Mpmos@6 vdd Q net@136 vdd PMOS L=0.6U W=3U AS=63.225P AD=13.95P PS=73.95U 
+PD=23.6U
Mpmos@7 vdd net@136 Q vdd PMOS L=0.6U W=3U AS=63.225P AD=13.95P PS=73.95U 
+PD=23.6U
Mpmos@8 vdd D net@221 vdd PMOS L=0.6U W=6U AS=7.425P AD=13.95P PS=12.3U 
+PD=23.6U
Mpmos@10 net@136 SAE B vdd PMOS L=0.6U W=67.5U AS=166.5P AD=63.225P PS=201.6U 
+PD=73.95U
Mpmos@11 Q SAE Bb vdd PMOS L=0.6U W=67.5U AS=144P AD=63.225P PS=171.6U 
+PD=73.95U
.ENDS SRAM_8x8__sense_amp

*** TOP LEVEL CELL: column4{lay}
Xcell2@0 net@246 net@260 gnd cell2@0_n cell2@0_q vdd net@479 Cell_Copy__cell2
Xcell2@7 net@246 net@260 gnd cell2@7_n cell2@7_q vdd net@254 Cell_Copy__cell2
Xcell2@8 net@246 net@260 gnd cell2@8_n cell2@8_q vdd net@268 Cell_Copy__cell2
Xcell2@9 net@246 net@260 gnd cell2@9_n cell2@9_q vdd net@271 Cell_Copy__cell2
Xcell2@10 net@246 net@260 gnd p40 o40 vdd net@281 Cell_Copy__cell2
Xcell2@11 net@246 net@260 gnd p50 o50 vdd net@290 Cell_Copy__cell2
Xcell2@12 net@246 net@260 gnd cell2@12_n cell2@12_q vdd net@298 
+Cell_Copy__cell2
Xcell2@13 net@246 net@260 gnd p70 o70 vdd net@302 Cell_Copy__cell2
Xcell2@14 net@355 net@365 gnd cell2@14_n cell2@14_q vdd net@479 
+Cell_Copy__cell2
Xcell2@15 net@355 net@365 gnd cell2@15_n cell2@15_q vdd net@254 
+Cell_Copy__cell2
Xcell2@16 net@355 net@365 gnd cell2@16_n cell2@16_q vdd net@268 
+Cell_Copy__cell2
Xcell2@17 net@355 net@365 gnd cell2@17_n cell2@17_q vdd net@271 
+Cell_Copy__cell2
Xcell2@18 net@355 net@365 gnd p41 cell2@18_q vdd net@281 Cell_Copy__cell2
Xcell2@19 net@355 net@365 gnd p51 cell2@19_q vdd net@290 Cell_Copy__cell2
Xcell2@20 net@355 net@365 gnd cell2@20_n cell2@20_q vdd net@298 
+Cell_Copy__cell2
Xcell2@21 net@355 net@365 gnd p71 cell2@21_q vdd net@302 Cell_Copy__cell2
Xcell2@22 net@791 net@792 gnd cell2@22_n cell2@22_q vdd net@479 
+Cell_Copy__cell2
Xcell2@23 net@791 net@792 gnd cell2@23_n cell2@23_q vdd net@254 
+Cell_Copy__cell2
Xcell2@24 net@791 net@792 gnd cell2@24_n cell2@24_q vdd net@268 
+Cell_Copy__cell2
Xcell2@25 net@791 net@792 gnd cell2@25_n cell2@25_q vdd net@271 
+Cell_Copy__cell2
Xcell2@26 net@791 net@792 gnd p42 cell2@26_q vdd net@281 Cell_Copy__cell2
Xcell2@27 net@791 net@792 gnd p52 cell2@27_q vdd net@290 Cell_Copy__cell2
Xcell2@28 net@791 net@792 gnd cell2@28_n cell2@28_q vdd net@298 
+Cell_Copy__cell2
Xcell2@29 net@791 net@792 gnd p72 cell2@29_q vdd net@302 Cell_Copy__cell2
Xcell2@30 net@901 net@917 gnd cell2@30_n cell2@30_q vdd net@479 
+Cell_Copy__cell2
Xcell2@31 net@901 net@917 gnd cell2@31_n cell2@31_q vdd net@254 
+Cell_Copy__cell2
Xcell2@32 net@901 net@917 gnd cell2@32_n cell2@32_q vdd net@268 
+Cell_Copy__cell2
Xcell2@33 net@901 net@917 gnd cell2@33_n cell2@33_q vdd net@271 
+Cell_Copy__cell2
Xcell2@34 net@901 net@917 gnd p43 cell2@34_q vdd net@281 Cell_Copy__cell2
Xcell2@35 net@901 net@917 gnd p53 cell2@35_q vdd net@290 Cell_Copy__cell2
Xcell2@36 net@901 net@917 gnd cell2@36_n cell2@36_q vdd net@298 
+Cell_Copy__cell2
Xcell2@37 net@901 net@917 gnd p73 cell2@37_q vdd net@302 Cell_Copy__cell2
Xcell2@38 net@981 net@980 gnd cell2@38_n cell2@38_q vdd net@479 
+Cell_Copy__cell2
Xcell2@39 net@981 net@980 gnd cell2@39_n cell2@39_q vdd net@254 
+Cell_Copy__cell2
Xcell2@40 net@981 net@980 gnd cell2@40_n cell2@40_q vdd net@268 
+Cell_Copy__cell2
Xcell2@41 net@981 net@980 gnd cell2@41_n cell2@41_q vdd net@271 
+Cell_Copy__cell2
Xcell2@42 net@981 net@980 gnd p44 cell2@42_q vdd net@281 Cell_Copy__cell2
Xcell2@43 net@981 net@980 gnd p54 cell2@43_q vdd net@290 Cell_Copy__cell2
Xcell2@44 net@981 net@980 gnd cell2@44_n cell2@44_q vdd net@298 
+Cell_Copy__cell2
Xcell2@45 net@981 net@980 gnd p74 cell2@45_q vdd net@302 Cell_Copy__cell2
Xcell2@46 net@1039 net@1037 gnd cell2@46_n cell2@46_q vdd net@479 
+Cell_Copy__cell2
Xcell2@47 net@1039 net@1037 gnd cell2@47_n cell2@47_q vdd net@254 
+Cell_Copy__cell2
Xcell2@48 net@1039 net@1037 gnd cell2@48_n cell2@48_q vdd net@268 
+Cell_Copy__cell2
Xcell2@49 net@1039 net@1037 gnd cell2@49_n cell2@49_q vdd net@271 
+Cell_Copy__cell2
Xcell2@50 net@1039 net@1037 gnd p45 cell2@50_q vdd net@281 Cell_Copy__cell2
Xcell2@51 net@1039 net@1037 gnd p55 cell2@51_q vdd net@290 Cell_Copy__cell2
Xcell2@52 net@1039 net@1037 gnd cell2@52_n cell2@52_q vdd net@298 
+Cell_Copy__cell2
Xcell2@53 net@1039 net@1037 gnd p75 cell2@53_q vdd net@302 Cell_Copy__cell2
Xcell2@54 net@1093 net@1094 gnd cell2@54_n cell2@54_q vdd net@479 
+Cell_Copy__cell2
Xcell2@55 net@1093 net@1094 gnd cell2@55_n cell2@55_q vdd net@254 
+Cell_Copy__cell2
Xcell2@56 net@1093 net@1094 gnd cell2@56_n cell2@56_q vdd net@268 
+Cell_Copy__cell2
Xcell2@57 net@1093 net@1094 gnd cell2@57_n cell2@57_q vdd net@271 
+Cell_Copy__cell2
Xcell2@58 net@1093 net@1094 gnd p46 cell2@58_q vdd net@281 Cell_Copy__cell2
Xcell2@59 net@1093 net@1094 gnd p56 cell2@59_q vdd net@290 Cell_Copy__cell2
Xcell2@60 net@1093 net@1094 gnd cell2@60_n cell2@60_q vdd net@298 
+Cell_Copy__cell2
Xcell2@61 net@1093 net@1094 gnd p76 cell2@61_q vdd net@302 Cell_Copy__cell2
Xcell2@62 net@1150 net@1149 gnd cell2@62_n cell2@62_q vdd net@479 
+Cell_Copy__cell2
Xcell2@63 net@1150 net@1149 gnd cell2@63_n cell2@63_q vdd net@254 
+Cell_Copy__cell2
Xcell2@64 net@1150 net@1149 gnd cell2@64_n cell2@64_q vdd net@268 
+Cell_Copy__cell2
Xcell2@65 net@1150 net@1149 gnd cell2@65_n cell2@65_q vdd net@271 
+Cell_Copy__cell2
Xcell2@66 net@1150 net@1149 gnd p47 o47 vdd net@281 Cell_Copy__cell2
Xcell2@67 net@1150 net@1149 gnd p57 o57 vdd net@290 Cell_Copy__cell2
Xcell2@68 net@1150 net@1149 gnd cell2@68_n cell2@68_q vdd net@298 
+Cell_Copy__cell2
Xcell2@69 net@1150 net@1149 gnd p77 o77 vdd net@302 Cell_Copy__cell2
Xdecoder@0 A B C DEN gnd net@7 net@6 net@5 net@4 net@3 net@2 net@1 net@0 vdd 
+SRAM_8x8__decoder
Xinv@0 gnd net@7 net@479 vdd inverter1__inv
Xinv@1 gnd net@6 net@254 vdd inverter1__inv
Xinv@2 gnd net@5 net@268 vdd inverter1__inv
Xinv@3 gnd net@4 net@271 vdd inverter1__inv
Xinv@4 gnd net@3 net@281 vdd inverter1__inv
Xinv@5 gnd net@2 net@290 vdd inverter1__inv
Xinv@6 gnd net@1 net@298 vdd inverter1__inv
Xinv@7 gnd net@0 net@302 vdd inverter1__inv
Mpmos@0 vdd P net@246 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@1 vdd P net@260 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@2 net@260 P net@246 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@24 vdd P net@355 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@25 vdd P net@365 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@26 net@365 P net@355 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@27 vdd P net@791 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@28 vdd P net@792 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@29 net@792 P net@791 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@30 vdd P net@901 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@31 vdd P net@917 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@32 net@917 P net@901 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@33 vdd P net@981 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@34 vdd P net@980 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@35 net@980 P net@981 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@36 vdd P net@1039 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@37 vdd P net@1037 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@38 net@1037 P net@1039 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@39 vdd P net@1093 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@40 vdd P net@1094 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@41 net@1094 P net@1093 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Mpmos@42 vdd P net@1150 vdd PMOS L=0.6U W=42U AS=38.992P AD=78.3P PS=86.85U 
+PD=118.8U
Mpmos@43 vdd P net@1149 vdd PMOS L=0.6U W=42U AS=58.05P AD=78.3P PS=88.8U 
+PD=118.8U
Mpmos@44 net@1149 P net@1150 vdd PMOS L=0.6U W=42U AS=38.992P AD=58.05P 
+PS=86.85U PD=88.8U
Xsense_am@0 net@246 net@260 d0 gnd q0 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@1 net@355 net@365 d1 gnd q1 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@2 net@791 net@792 d2 gnd q2 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@3 net@901 net@917 d3 gnd q3 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@4 net@981 net@980 d4 gnd q4 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@5 net@1039 net@1037 d5 gnd q5 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@6 net@1093 net@1094 d6 gnd q6 SAE vdd WE SRAM_8x8__sense_amp
Xsense_am@7 net@1150 net@1149 d7 gnd q7 SAE vdd WE SRAM_8x8__sense_amp

* Spice Code nodes in cell cell 'column4{lay}'
vdd vdd 0 dc 5
va A 0 DC 0 pwl 100n 0 110n 5 150n 5 160n 0 200n 0 210n 5
vb B 0 DC 0 pwl 100n 5 110n 0 200n 0 210n 5 350n 5 360n 0 500n 0 510n 5
vc C 0 DC 0 pwl 100n 0 110n 5 350n 5 360n 0 500n 0 510n 5
vp P 0 DC 0 pwl 50n 5 60n 0 100n 0 110n 5 200n 5 210n 0 250n 0 260n 5 350n 5 
+360n 0 400n 0 410n 5 500n 5 510n 0 550n 0 560n 5
vwe WE 0 DC 0 pwl 100n 5 110n 0 250n 0 260n 5 300n 5 310n 0
vsae SAE 0 DC 0 pwl 100n 5 110n 0 150n 0 160n 5 250n 5 260n 0 300n 0 310n 5 
+400n 5 410n 0 450n 0 460n 5 550n 5 560n 0 600n 0 610n 5
vden DEN 0 dc 0 pwl 100n 0 110n 5 150n 5 160n 0 250n 0 260n 5 300n 5 310n 0 
+400n 0 410n 5 450n 5 460n 0 550n 0 560n 5 600n 5 610n 0
vd0 d0 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd1 d1 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd2 d2 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd3 d3 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd4 d4 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd5 d5 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd6 d6 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
vd7 d7 0 dc 0 pwl 200n 0 210n 5 300n 5 310n 0
.IC V(p50)=0 V(p51)=0 V(p52)=0 V(p53)=0 V(p54)=0 V(p55)=0 V(p56)=0 V(p57)=0 
+V(p40)=0 V(p41)=0 V(p42)=0 V(p43)=0 V(p44)=0 V(p45)=0 V(p46)=0 V(p47)=0 
+V(p70)=0 V(p71)=0 V(p72)=0 V(p73)=0 V(p74)=0 V(p75)=0 V(p76)=0 V(p77)=0
.tran 0 800ns
.include C5_models.txt
.END
